library verilog;
use verilog.vl_types.all;
entity NanoControlador_vlg_vec_tst is
end NanoControlador_vlg_vec_tst;
