library verilog;
use verilog.vl_types.all;
entity port_and_vlg_vec_tst is
end port_and_vlg_vec_tst;
