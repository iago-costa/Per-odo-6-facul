library ieee; --DEFINICAO DA BIBLIOTECA IEEE para usar definicoes do tipo bit booleano entre outras coisas
USE ieee.std_logic_1164.all; --DECLARACAO NECESSARIA PARA USAR OS DADOS CORRESPONDENTES A LÓGICA PADRAO DA BIBLIOTECA
ENTITY dff_logic IS --DECLARACAO DA ENTIDADE CONTENDO OS PINOS I/0.
PORT (d,clk:IN BIT; --DECLARACAO DAS ENTRADAS D E CLOCK DE TIPOS BITS
		q:OUT BIT); --DECLARACAO DA SAIDA Q DO TIPO BIT
END dff_logic; -- FIM DA DEFINICAO DA ENTIDADE
ARCHITECTURE behavior OF dff_logic IS --DECLARACAO DA ARQUITEUTURA, OU SEJA, A LÓGICA DO CIRCUITO
BEGIN  --INICIO DA ARQUITETURA
	PROCESS(clk) --CLK CORRESPONDE A LISTA DE SINAIS QUE PODEM ALTERAR A SAIDA DO CIRCUITO
	BEGIN --Inicio da descricao logica do processo
		IF(clk'event AND clk = '1') THEN	--INICIO DA CONDICIONAL
		q <= d; --ACAO QUE DEVERA FAZER CASO A CONDICAO SEJA FAVORECIDA
		END IF; --FIM DA CONDICIONAL
	END PROCESS; --FIM DO PROCESSO
END behavior; --FIM DA ARQUITETURA, OU SEJA, DA LÓGICA DO CIRCUITO
		