library verilog;
use verilog.vl_types.all;
entity dff_logic_reset_vlg_vec_tst is
end dff_logic_reset_vlg_vec_tst;
